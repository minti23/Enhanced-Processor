LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY DFFp IS 
PORT ( CLK: IN STD_LOGIC;
		 D: IN STD_LOGIC;
		 Q: OUT STD_LOGIC;
		 RESET: IN STD_LOGIC;
		 EN: IN STD_LOGIC);
END ENTITY;

ARCHITECTURE BEH OF DFFp IS

BEGIN
	PROCESS (CLK, RESET, EN)
	BEGIN
	IF rising_edge(CLK) AND (EN ='1') THEN
	Q <= D;
	END IF;
	IF RESET ='1' THEN
	Q <= '0';
	END IF;
	END PROCESS;
END BEH;